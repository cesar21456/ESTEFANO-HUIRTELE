module PC(input clk,input[31:0] pc,output[31:0] direccion);

assign direccion=pc;
endmodule

